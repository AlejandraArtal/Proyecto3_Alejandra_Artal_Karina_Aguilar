`timescale 1ns / 1ps

module font_rom_caracteres
(
    input wire [10:0] addr,
    output reg [15:0] data = 16'd0
);

always @ * begin
    data = 16'd0;
    case (addr)
	 //code x00
      11'h0: data = 16'b0000000000000000;
      11'h1: data = 16'b0000000000000000;
      11'h2: data = 16'b0000000000000000;
      11'h3: data = 16'b0000000000000000;
      11'h4: data =  16'b0000000000000000;
      11'h5: data =  16'b0000000000000000;
      11'h6: data =  16'b0000000000000000;
      11'h7: data =  16'b0000000000000000;
      11'h8: data =  16'b0000000000000000;
      11'h9: data =  16'b0000011111110000;
      11'ha: data =  16'b0000111111111100;
      11'hb: data =  16'b0001111111111110;
      11'hc: data =  16'b0011111111111110;
      11'hd: data =  16'b0111111111111111;
      11'he: data =  16'b0111111100111111;
      11'hf: data =  16'b0111111000011111;
      11'h10: data = 16'b0111111000011111;
      11'h11: data = 16'b0111111000011111;
      11'h12: data = 16'b0111111100111111;
      11'h13: data = 16'b0111111111111111;
      11'h14: data = 16'b0011111111111110;
      11'h15: data = 16'b0001111111111110;
      11'h16: data = 16'b0000111111111100;
      11'h17: data = 16'b0000011111110000;
      11'h18: data = 16'b0000000000000000;
      11'h19: data = 16'b0000000000000000;
      11'h1a: data = 16'b0000000000000000;
      11'h1b: data = 16'b0000000000000000;
      11'h1c: data = 16'b0000000000000000;
      11'h1d: data = 16'b0000000000000000;
      11'h1e: data = 16'b0000000000000000;
      11'h1f: data = 16'b0000000000000000;
		
		//code x01
      11'h20: data = 16'b0000000000000000;
      11'h21: data = 16'b0000000000000000;
      11'h22: data = 16'b0000000000000000;
      11'h23: data = 16'b0000000000000000;
      11'h24: data = 16'b0000000000000000;
      11'h25: data = 16'b0000000000000000;
      11'h26: data = 16'b0000000000000000;
      11'h27: data = 16'b0000000000000000;
      11'h28: data = 16'b0000000000000000;
      11'h29: data = 16'b0000000111100000;
      11'h2a: data = 16'b0000001111100000;
      11'h2b: data = 16'b0000111111100000;
      11'h2c: data = 16'b0000111111100000;
      11'h2d: data = 16'b0000111111100000;
      11'h2e: data = 16'b0000111111100000;
      11'h2f: data = 16'b0000111111100000;
      11'h30: data = 16'b0000001111100000;
      11'h31: data = 16'b0000001111100000;
      11'h32: data = 16'b0000001111100000;
      11'h33: data = 16'b0000001111100000;
      11'h34: data = 16'b0000001111100000;
      11'h35: data = 16'b0000001111100000;
      11'h36: data = 16'b0000001111100000;
      11'h37: data = 16'b0000001111100000;
      11'h38: data = 16'b0000000000000000;
      11'h39: data = 16'b0000000000000000;
      11'h3a: data = 16'b0000000000000000;
      11'h3b: data = 16'b0000000000000000;
      11'h3c: data = 16'b0000000000000000;
      11'h3d: data = 16'b0000000000000000;
      11'h3e: data = 16'b0000000000000000;
      11'h3f: data = 16'b0000000000000000;
		
		//code x02
		11'h40: data = 16'b0000000000000000;
      11'h41: data = 16'b0000000000000000;
      11'h42: data = 16'b0000000000000000;
      11'h43: data = 16'b0000000000000000;
      11'h44: data = 16'b0000000000000000;
      11'h45: data = 16'b0000000000000000;
      11'h46: data = 16'b0000000000000000;
      11'h47: data = 16'b0000000000000000;
      11'h48: data = 16'b0000000000000000;
      11'h49: data = 16'b0000111111110000;
      11'h4a: data = 16'b0011111111111000;
      11'h4b: data = 16'b0011111111111100;
      11'h4c: data = 16'b0011111111111100;
      11'h4d: data = 16'b0011110011111100;
      11'h4e: data = 16'b0000000001111100;
      11'h4f: data = 16'b0000000001111100;
      11'h50: data = 16'b0000000011111000;
      11'h51: data = 16'b0000000111110000;
      11'h52: data = 16'b0000001111100000;
      11'h53: data = 16'b0000111111000000;
      11'h54: data = 16'b0011111111111110;
      11'h55: data = 16'b0011111111111110;
      11'h56: data = 16'b0011111111111110;
      11'h57: data = 16'b0011111111111110;
      11'h58: data = 16'b0000000000000000;
      11'h59: data = 16'b0000000000000000;
      11'h5a: data = 16'b0000000000000000;
      11'h5b: data = 16'b0000000000000000;
      11'h5c: data = 16'b0000000000000000;
      11'h5d: data = 16'b0000000000000000;
      11'h5e: data = 16'b0000000000000000;
      11'h5f: data = 16'b0000000000000000;
		
		//code x03
		11'h60: data = 16'b0000000000000000;
      11'h61: data = 16'b0000000000000000;
      11'h62: data = 16'b0000000000000000;
      11'h63: data = 16'b0000000000000000;
      11'h64: data = 16'b0000000000000000;
      11'h65: data = 16'b0000000000000000;
      11'h66: data = 16'b0000000000000000;
      11'h67: data = 16'b0000000000000000;
      11'h68: data = 16'b0000000000000000;
      11'h69: data = 16'b0001111111110000;
      11'h6a: data = 16'b0001111111111000;
      11'h6b: data = 16'b0001111111111000;
      11'h6c: data = 16'b0001111111111000;
      11'h6d: data = 16'b0000000111111000;
      11'h6e: data = 16'b0000111111111000;
      11'h6f: data = 16'b0000111111110000;
      11'h70: data = 16'b0000111111111000;
      11'h71: data = 16'b0000000011111100;
      11'h72: data = 16'b0000000011111100;
      11'h73: data = 16'b0001110011111100;
      11'h74: data = 16'b0011111111111100;
      11'h75: data = 16'b0011111111111100;
      11'h76: data = 16'b0011111111111000;
      11'h77: data = 16'b0001111111110000;
      11'h78: data = 16'b0000000000000000;
      11'h79: data = 16'b0000000000000000;
      11'h7a: data = 16'b0000000000000000;
      11'h7b: data = 16'b0000000000000000;
      11'h7c: data = 16'b0000000000000000;
      11'h7d: data = 16'b0000000000000000;
      11'h7e: data = 16'b0000000000000000;
      11'h7f: data = 16'b0000000000000000;
		
		//code x04
		11'h80: data = 16'b0000000000000000;
      11'h81: data = 16'b0000000000000000;
      11'h82: data = 16'b0000000000000000;
      11'h83: data = 16'b0000000000000000;
      11'h84: data = 16'b0000000000000000;
      11'h85: data = 16'b0000000000000000;
      11'h86: data = 16'b0000000000000000;
      11'h87: data = 16'b0000000000000000;
      11'h88: data = 16'b0000000000000000;
      11'h89: data = 16'b0000000111111000;
      11'h8a: data = 16'b0000001111111000;
      11'h8b: data = 16'b0000001111111000;
      11'h8c: data = 16'b0000011111111000;
      11'h8d: data = 16'b0000111111111000;
      11'h8e: data = 16'b0000111111111000;
      11'h8f: data = 16'b0001111011111000;
      11'h90: data = 16'b0011111011111000;
      11'h91: data = 16'b0111110011111000;
      11'h92: data = 16'b0111111111111100;
      11'h93: data = 16'b0111111111111100;
      11'h94: data = 16'b0111111111111100;
      11'h95: data = 16'b0000000111111000;
      11'h96: data = 16'b0000000111111000;
      11'h97: data = 16'b0000000111111000;
      11'h98: data = 16'b0000000000000000;
      11'h99: data = 16'b0000000000000000;
      11'h9a: data = 16'b0000000000000000;
      11'h9b: data = 16'b0000000000000000;
      11'h9c: data = 16'b0000000000000000;
      11'h9d: data = 16'b0000000000000000;
      11'h9e: data = 16'b0000000000000000;
      11'h9f: data = 16'b0000000000000000;
		
		//code x05
		11'ha0: data = 16'b0000000000000000;
      11'ha1: data = 16'b0000000000000000;
      11'ha2: data = 16'b0000000000000000;
      11'ha3: data = 16'b0000000000000000;
      11'ha4: data = 16'b0000000000000000;
      11'ha5: data = 16'b0000000000000000;
      11'ha6: data = 16'b0000000000000000;
      11'ha7: data = 16'b0000000000000000;
      11'ha8: data = 16'b0000000000000000;
      11'ha9: data = 16'b0001111111111000;
      11'haa: data = 16'b0001111111111000;
      11'hab: data = 16'b0001111111111000;
      11'hac: data = 16'b0001111111110000;
      11'had: data = 16'b0001111000000000;
      11'hae: data = 16'b0001111111110000;
      11'haf: data = 16'b0001111111111000;
      11'hb0: data = 16'b0001111111111100;
      11'hb1: data = 16'b0000000011111100;
      11'hb2: data = 16'b0000000001111100;
      11'hb3: data = 16'b0000000011111100;
      11'hb4: data = 16'b0011111111111100;
      11'hb5: data = 16'b0011111111111100;
      11'hb6: data = 16'b0011111111111000;
      11'hb7: data = 16'b0011111111110000;
      11'hb8: data = 16'b0000000000000000;
      11'hb9: data = 16'b0000000000000000;
      11'hba: data = 16'b0000000000000000;
      11'hbb: data = 16'b0000000000000000;
      11'hbc: data = 16'b0000000000000000;
      11'hbd: data = 16'b0000000000000000;
      11'hbe: data = 16'b0000000000000000;
      11'hbf: data = 16'b0000000000000000;
		
		//code x06
		11'hc0: data = 16'b0000000000000000;
      11'hc1: data = 16'b0000000000000000;
      11'hc2: data = 16'b0000000000000000;
      11'hc3: data = 16'b0000000000000000;
      11'hc4: data = 16'b0000000000000000;
      11'hc5: data = 16'b0000000000000000;
      11'hc6: data = 16'b0000000000000000;
      11'hc7: data = 16'b0000000000000000;
      11'hc8: data = 16'b0000000000000000;
      11'hca: data = 16'b0000111111111100;
      11'hcb: data = 16'b0011111111111110;
      11'hcc: data = 16'b0011111111111110;
      11'hcd: data = 16'b0011111100000000;
      11'hce: data = 16'b0011111011111000;
      11'hcf: data = 16'b0011111111111100;
      11'hd0: data = 16'b0011111111111100;
      11'hd1: data = 16'b0011111001111110;
      11'hd2: data = 16'b0011111000111110;
      11'hd3: data = 16'b0011111001111110;
      11'hd4: data = 16'b0011111111111110;
      11'hd5: data = 16'b0011111111111110;
      11'hd6: data = 16'b0011111111111110;
      11'hd7: data = 16'b0001111111111100;
      11'hd8: data = 16'b0000000000000000;
      11'hd9: data = 16'b0000000000000000;
      11'hda: data = 16'b0000000000000000;
      11'hdb: data = 16'b0000000000000000;
      11'hdc: data = 16'b0000000000000000;
      11'hdd: data = 16'b0000000000000000;
      11'hde: data = 16'b0000000000000000;
      11'hdf: data = 16'b0000000000000000;
		
		//code x07
		11'he0: data = 16'b0000000000000000;
      11'he1: data = 16'b0000000000000000;
      11'he2: data = 16'b0000000000000000;
      11'he3: data = 16'b0000000000000000;
      11'he4: data = 16'b0000000000000000;
      11'he5: data = 16'b0000000000000000;
      11'he6: data = 16'b0000000000000000;
      11'he7: data = 16'b0000000000000000;
      11'he8: data = 16'b0000000000000000;
      11'he9: data = 16'b0011111111111100;
      11'hea: data = 16'b0011111111111100;
      11'heb: data = 16'b0011111111111100;
      11'hec: data = 16'b0011111111111100;
      11'hed: data = 16'b0000000111111000;
      11'hee: data = 16'b0000000111110000;
      11'hef: data = 16'b0000001111110000;
      11'hf0: data = 16'b0000001111100000;
      11'hf1: data = 16'b0000011111100000;
      11'hf2: data = 16'b0000011111000000;
      11'hf3: data = 16'b0000011111000000;
      11'hf4: data = 16'b0000111111000000;
      11'hf5: data = 16'b0000111111000000;
      11'hf6: data = 16'b0000111111000000;
      11'hf7: data = 16'b0000111111000000;
      11'hf8: data = 16'b0000000000000000;
      11'hf9: data = 16'b0000000000000000;
      11'hfa: data = 16'b0000000000000000;
      11'hfb: data = 16'b0000000000000000;
      11'hfc: data = 16'b0000000000000000;
      11'hfd: data = 16'b0000000000000000;
      11'hfe: data = 16'b0000000000000000;
      11'hff: data = 16'b0000000000000000;
		
		//code x08
		11'h100: data = 16'b0000000000000000;
      11'h101: data = 16'b0000000000000000;
      11'h102: data = 16'b0000000000000000;
      11'h103: data = 16'b0000000000000000;
      11'h104: data = 16'b0000000000000000;
      11'h105: data = 16'b0000000000000000;
      11'h106: data = 16'b0000000000000000;
      11'h107: data = 16'b0000000000000000;
      11'h108: data = 16'b0000000000000000;
      11'h109: data = 16'b0000111111110000;
      11'h10a: data = 16'b0001111111111000;
      11'h10b: data = 16'b0001111111111100;
      11'h10c: data = 16'b0011111001111100;
      11'h10d: data = 16'b0011111000111100;
      11'h10e: data = 16'b0011111100111100;
      11'h10f: data = 16'b0001111111111000;
      11'h110: data = 16'b0001111111111000;
      11'h111: data = 16'b0001111111111100;
      11'h112: data = 16'b0011110011111100;
      11'h113: data = 16'b0011110000111100;
      11'h114: data = 16'b0011111001111100;
      11'h115: data = 16'b0011111111111100;
      11'h116: data = 16'b0001111111111000;
      11'h117: data = 16'b0000111111110000;
      11'h118: data = 16'b0000000000000000;
      11'h119: data = 16'b0000000000000000;
      11'h11a: data = 16'b0000000000000000;
      11'h11b: data = 16'b0000000000000000;
      11'h11c: data = 16'b0000000000000000;
      11'h11d: data = 16'b0000000000000000;
      11'h11e: data = 16'b0000000000000000;
      11'h11f: data = 16'b0000000000000000;
		
		//code x09
		11'h120: data = 16'b0000000000000000;
      11'h121: data = 16'b0000000000000000;
      11'h122: data = 16'b0000000000000000;
      11'h123: data = 16'b0000000000000000;
      11'h124: data = 16'b0000000000000000;
      11'h125: data = 16'b0000000000000000;
      11'h126: data = 16'b0000000000000000;
      11'h127: data = 16'b0000000000000000;
      11'h128: data = 16'b0000000000000000;
      11'h129: data = 16'b0000111111110000;
      11'h12a: data = 16'b0001111111111000;
      11'h12b: data = 16'b0011111111111100;
      11'h12c: data = 16'b0111111111111100;
      11'h12d: data = 16'b0111110001111110;
      11'h12e: data = 16'b0111100000111111;
      11'h12f: data = 16'b0111110001111111;
      11'h130: data = 16'b0011111111111110;
      11'h131: data = 16'b0011111111111100;
      11'h132: data = 16'b0001111111111100;
      11'h133: data = 16'b0000111111111100;
      11'h134: data = 16'b0000011111111000;
      11'h135: data = 16'b0011111111110000;
      11'h136: data = 16'b0011111111100000;
      11'h137: data = 16'b0001111110000000;
      11'h138: data = 16'b0000000000000000;
      11'h139: data = 16'b0000000000000000;
      11'h13a: data = 16'b0000000000000000;
      11'h13b: data = 16'b0000000000000000;
      11'h13c: data = 16'b0000000000000000;
      11'h13d: data = 16'b0000000000000000;
      11'h13e: data = 16'b0000000000000000;
      11'h13f: data = 16'b0000000000000000;
		
		//code x10
		11'h140: data = 16'b0000000000000000;
      11'h141: data = 16'b0000000000000000;
      11'h142: data = 16'b0000000000000000;
      11'h143: data = 16'b0000000000000000;
      11'h144: data = 16'b0000000000000000;
      11'h145: data = 16'b0000000000000000;
      11'h146: data = 16'b0000000000000000;
      11'h147: data = 16'b0000000000000000;
      11'h148: data = 16'b0000000000000000;
      11'h149: data = 16'b0000000000000000;
      11'h14a: data = 16'b0000000000000000;
      11'h14b: data = 16'b0000001111000000;
      11'h14c: data = 16'b0000001111100000;
      11'h14d: data = 16'b0000011111100000;
      11'h14e: data = 16'b0000001111100000;
      11'h14f: data = 16'b0000001111000000;
      11'h150: data = 16'b0000000000000000;
      11'h151: data = 16'b0000001111000000;
      11'h152: data = 16'b0000001111100000;
      11'h153: data = 16'b0000011111100000;
      11'h154: data = 16'b0000001111100000;
      11'h155: data = 16'b0000001111000000;
      11'h156: data = 16'b0000000000000000;
      11'h157: data = 16'b0000000000000000;
      11'h158: data = 16'b0000000000000000;
      11'h159: data = 16'b0000000000000000;
      11'h15a: data = 16'b0000000000000000;
      11'h15b: data = 16'b0000000000000000;
      11'h15c: data = 16'b0000000000000000;
      11'h15d: data = 16'b0000000000000000;
      11'h15e: data = 16'b0000000000000000;
      11'h15f: data = 16'b0000000000000000;
		
		//code x11
		11'h160: data = 16'b0000000000000000;
      11'h161: data = 16'b0000000000000000;
      11'h162: data = 16'b0000000000000000;
      11'h163: data = 16'b0000000000000000;
      11'h164: data = 16'b0000000000000000;
      11'h165: data = 16'b0000000000000000;
      11'h166: data = 16'b0000000000000000;
      11'h167: data = 16'b0000000000000000;
		11'h168: data = 16'b0000000000000000;
      11'h169: data = 16'b0000000000000000;
      11'h16a: data = 16'b0000000000000000;
      11'h16b: data = 16'b0000000000000000;
      11'h16c: data = 16'b0000000000000000;
      11'h16d: data = 16'b0000000000000000;
      11'h16e: data = 16'b0000000000000000;
      11'h16f: data = 16'b0000000000000000;
		11'h170: data = 16'b0000000000000000;
      11'h171: data = 16'b0000000000000000;
      11'h172: data = 16'b0000000000000000;
      11'h173: data = 16'b0000000000000000;
      11'h174: data = 16'b0000000000000000;
      11'h175: data = 16'b0000000000000000;
      11'h176: data = 16'b0000000000000000;
      11'h177: data = 16'b0000000000000000;
		11'h178: data = 16'b0000000000000000;
      11'h179: data = 16'b0000000000000000;
		11'h17a: data = 16'b0000000000000000;
      11'h17b: data = 16'b0000000000000000;
      11'h17c: data = 16'b0000000000000000;
      11'h17d: data = 16'b0000000000000000;
      11'h17e: data = 16'b0000000000000000;
      11'h17f: data = 16'b0000000000000000;
		
		endcase
end

endmodule
